package game_constants_pkg;
  parameter int POSITION_CHANGE_FREQ_IN_CLOCKS = 10;
  parameter int DEBOUNCE_WIDTH_IN_CLOCKS       = 8;
  parameter int TOTAL_WIDTH                    = 640;
  parameter int TOTAL_HEIGHT                   = 480;
  parameter int PADDLE_DISTANCE_FROM_EDGE      = 40;
  parameter int PADDLE_HEIGHT                  = 100;
  parameter int PADDLE_WIDTH                   = 15;
  parameter int BALL_SIDE_SIZE                 = 24;
endpackage